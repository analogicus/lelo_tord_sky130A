*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_dac_lpe.spi
#else
.include ../../../work/xsch/TB_dac.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

.param f_CLK = 1MegHz
.param T_CLK = {1/f_CLK}

.param TD = {T_CLK*3}
.param TR = {T_CLK/100}
.param TF = {TR}
.param PW = {T_CLK}
.param PER = {T_CLK}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0    DC 0
VDD  VDD  VSS  DC {AVDD}
VSLP SLP  VSS  PWL 0.25us {AVDD} 0.3us 0V

VB0  B0   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*8/16} {PER})
VB1  B1   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*9/16} {PER})
VB2  B2   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*10/16} {PER})
VB3  B3   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*11/16} {PER})
VB4  B4   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*12/16} {PER})
VB5  B5   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*13/16} {PER})
VB6  B6   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*14/16} {PER})
VB7  B7   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*15/16} {PER})

VBT  BT   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*8/16} {PER})
* VBT  BT   VSS  DC 0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
* .include ../svinst.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

echo "T_CLK = " {T_CLK}


optran 0 0 0 1n 1u 0


tran 1n 15us 1p
write
quit


.endc

.end
