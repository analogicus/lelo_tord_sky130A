*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/dig-to-time_lpe.spi
#else
.include ../../../work/xsch/dig-to-time.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param f_CLK = 1MegHz
.param T_CLK = {1/f_CLK}
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0    dc 0
VDD  VDD  VSS  pwl 0 0 10n {AVDD}
VRST RST  VSS  pwl 1.3us {AVDD} 1.9us 0V 
VCLK CLK  VSS  pulse(0V {AVDD} {T_CLK/10} {T_CLK/100} {T_CLK/100} {T_CLK/2} {T_CLK})

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names
VB0 d.0 d0 dc 0
VB1 d.1 d1 dc 0
VB2 d.2 d2 dc 0
VB3 d.3 d3 dc 0

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.option savecurrents
.save all

.save v(vdd) v(vss)
.save v(clk) v(rst)
.save v(d0) v(d1) v(d2) v(d3)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

optran 0 0 0 1n 1u 0


tran 1n 20us 1p
write
quit


.endc

.end
