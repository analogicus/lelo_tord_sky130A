*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_gm_lpe.spi
#else
.include ../../../work/xsch/TB_gm.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VGND VD 0   dc 0
VSG VS  VG  dc 1.0V
VSD VS  VD  dc 1.8V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.option savecurrents
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


op

dc VSG 0 1.8 0.01

set fend = .out
set wr_singlescale
set wr_vecnames
option numdgt = 5
echo writing to {cicname}{$fend}

wrdata {cicname}{$fend}
+ v(vs) v(vg) v(vd)
+ i(v.xdut.v1) i(v.xdut.v2) i(v.xdut.v3) i(v.xdut.v4)
* + i(vs) i(vg) i(vd)
 

quit

.endc

.end
