magic
tech sky130A
timestamp 1770504968
<< locali >>
rect 2744 2544 2840 2584
<< metal1 >>
rect 2036 5164 2132 5204
rect 2228 4084 2324 4124
rect 6728 4084 6824 4124
rect 2872 2544 2904 2584
rect 5572 2544 5604 2584
use cmp_two_stage_nmos_cross_coupled  x1 ../LELO_TORD_SKY130A
timestamp 1770504890
transform 1 0 0 0 1 0
box -200 -13 7060 5800
<< labels >>
flabel locali s 2744 2544 2840 2584 0 FreeSans 200 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal1 s 2036 5164 2132 5204 0 FreeSans 200 0 0 0 VDD
port 2 nsew power bidirectional
flabel metal1 s 2872 2544 2904 2584 0 FreeSans 200 0 0 0 VIN
port 3 nsew signal bidirectional
flabel metal1 s 5572 2544 5604 2584 0 FreeSans 200 0 0 0 VIP
port 4 nsew signal bidirectional
flabel metal1 s 6728 4084 6824 4124 0 FreeSans 200 0 0 0 VOUT
port 5 nsew signal bidirectional
flabel metal1 s 2228 4084 2324 4124 0 FreeSans 200 0 0 0 VOUT_N
port 6 nsew signal bidirectional
flabel space 3584 3638 3612 3671 0 FreeSans 800 0 0 0 VIPDRN
port 7 nsew
flabel space 5324 3642 5352 3675 0 FreeSans 800 0 0 0 VINDRN
port 8 nsew
flabel space 4395 2116 4423 2149 0 FreeSans 800 0 0 0 VSRC
port 9 nsew
flabel space 684 3397 712 3430 0 FreeSans 800 0 0 0 VBIAS
<< properties >>
string FIXED_BBOX 0 0 6824 8000
<< end >>
