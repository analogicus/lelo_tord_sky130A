*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bgr_core_lpe.spi
#else
.include ../../../work/xsch/bgr_core.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3
* .option method=gear

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD    VDD       VSS DC  {AVDD}
VCTRL  CTRL      VSS PWL 0ns 0V 10ns {AVDD}
VSW1   SWBRANCH1 VSS PULSE(0V {AVDD} 1ns 1ps 1ps 999ps 2ns)
VSW2   SWBRANCH2 VSS PULSE({AVDD} 0V 1ns 1ps 1ps 999ps 2ns)
VCAP1  SWCAP1    VSS DC  {AVDD}
VCAP2  SWCAP2    VSS DC  {AVDD}
VREF1  SWREF1    VSS DC  0V
VREF2  SWREF2    VSS DC  0V
VDRAIN SWDRAIN   VSS PWL 0ns {AVDD} 900ps 0V
VSS    VSS       0   DC  0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.options savecurrents
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1ns 10ns 1ps
write
quit


.endc

.end
