*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_dac_lpe.spi
#else
.include ../../../work/xsch/TB_dac.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param f_CLK = 32MegHz
.param T_CLK = {1/f_CLK}

.param AVDD = {vdda}

.param f_CLK2 = 200kHz
.param T_CLK2 = {1/f_CLK2}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0 dc 0
VDD VDD VSS dc {AVDD}

VD0 d0 vss dc 0V
VD1 d1 vss dc 0V
VD2 d2 vss dc 0V
VD3 d3 vss pwl 100ns 0V 100.1ns {AVDD}
VCLK CLK VSS pulse(0V {AVDD} {T_CLK/10} {T_CLK/10000} {T_CLK/10000} {T_CLK/2} {T_CLK})

VDACCLK dac_CLK VSS pulse(0V {AVDD} {T_CLK2/10} {T_CLK2/100} {T_CLK2/100} {T_CLK2/2} {T_CLK2})
VRST dac_RST VSS pwl 1.3us {AVDD} 1.9us 0V 
VSLEEP SLEEP VSS pwl 0.25us {AVDD} 0.3us 0V


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names

VB0 b.0 b0 dc 0
VB1 b.1 b1 dc 0
VB2 b.2 b2 dc 0
VB3 b.3 b3 dc 0

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
*.option savecurrents

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

* Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

optran 0 0 0 1n 1u 0


tran 1n 75us 1p
write
quit


.endc

.end
