*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_temp_sens_lpe.spi
#else
.include ../../../work/xsch/TB_temp_sens.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10ps
.param AVDD = {vdda}

.csparam voltage_supply = {vdda}

* Circuit temperature given in degrees Celsius
.csparam circuit_temperature = -40
.param finetuning_frequency = 2
.param dutycycle = 55

* Finetuning frequency given in Mega Hertz and periode given in micro seconds
.csparam clock_frequency = {finetuning_frequency}
.csparam clock_periode = {1/finetuning_frequency}

* clock_frequency = 2 MHz => clock_periode = 0.5 us
* clock_frequency = 1 MHz => clock_periode = 1.0 us
.param f_clk = {finetuning_frequency * 1MegHz}
.param T_clk = {1/f_clk}
.param TD = {T_clk}
.param TR = {T_clk/100}
.param TF = {TR}
.param PW = {T_clk}
.param PER = {T_clk}

* Time averaging duty cycle is given in percent
.param ratio = {dutycycle/100}
.csparam duty_cycle = {dutycycle}

* Stepping Current out of DAC
.param step_start = 6.0us
.param step_length = {4*T_clk}
.csparam simulation_length = {step_start + 5*step_length}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS   VSS   0    dc 0V
VDD   VDD   VSS  dc {AVDD}
VSLP  SLP VSS pwl 0.02us {AVDD} 0.03us 0V

* VB0  B0   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*8/16} {PER})
* VB1  B1   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*9/16} {PER})
* VB2  B2   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*10/16} {PER})
* VB3  B3   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*11/16} {PER})
* VB4  B4   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*12/16} {PER})
* VB5  B5   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*13/16} {PER})
* VB6  B6   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*14/16} {PER})
* VB7  B7   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*15/16} {PER})

VB0  B0   VSS  dc pwl {step_start + 0*step_length} 0V {step_start + 0*step_length + 0.01us} {AVDD}
VB1  B1   VSS  dc pwl {step_start + 1*step_length} 0V {step_start + 1*step_length + 0.01us} {AVDD}
VB2  B2   VSS  dc pwl {step_start + 2*step_length} 0V {step_start + 2*step_length + 0.01us} {AVDD}
VB3  B3   VSS  dc pwl {step_start + 3*step_length} 0V {step_start + 3*step_length + 0.01us} {AVDD}
VB4  B4   VSS  dc pwl {step_start + 4*step_length} 0V {step_start + 4*step_length + 0.01us} {AVDD}
* VB5  B5   VSS  dc pwl {step_start + 5*step_length} 0V {step_start + 5*step_length + 0.01us} {AVDD}
* VB6  B6   VSS  dc pwl {step_start + 6*step_length} 0V {step_start + 6*step_length + 0.01us} {AVDD}
* VB7  B7   VSS  dc pwl {step_start + 7*step_length} 0V {step_start + 7*step_length + 0.01us} {AVDD}

* VB0  B0   VSS  dc 0V
* VB1  B1   VSS  dc 0V
* VB2  B2   VSS  dc 0V
* VB3  B3   VSS  dc 0V
* VB4  B4   VSS  dc 0V
VB5  B5   VSS  dc 0V
VB6  B6   VSS  dc 0V
VB7  B7   VSS  dc 0V

* VBT  BT   VSS  PULSE({AVDD} 0V {2*TD} {TR} {TF} {PW*ratio} {PER})
VBT  BT   VSS  PULSE(0V {AVDD} {2*TD} {TR} {TF} {PW*ratio} {PER})
* VBT  BT   VSS  DC 0V

VSWBRANCH1 SWBRN1 VSS dc {AVDD}
VSWBRANCH2 SWBRN2 VSS dc {AVDD}
VSWBRANCH3 SWBRN3 VSS dc {AVDD}
* VSWBRANCH1 SWBRN1 VSS dc 0
* VSWBRANCH2 SWBRN2 VSS dc 0
* VSWBRANCH3 SWBRN3 VSS dc 0

* VSWBGR1 SWBGR1 VSS dc {AVDD}
* VSWBGR2 SWBGR2 VSS dc {AVDD}
VSWBGR1 SWBGR1 VSS dc 0
VSWBGR2 SWBGR2 VSS dc 0

* VSWCAP1 SWCAP1 VSS dc {AVDD}
* VSWCAP2 SWCAP2 VSS dc {AVDD}
* VSWCAP3 SWCAP3 VSS dc {AVDD}
* VSWCAP1 SWCAP1 VSS dc 0
* VSWCAP2 SWCAP2 VSS dc 0
* VSWCAP3 SWCAP3 VSS dc 0
VSWCAP1 SWCAP1 VSS pwl 0.09us 0V 0.1us {AVDD} 
VSWCAP2 SWCAP2 VSS pwl 0.09us 0V 0.1us {AVDD} 
VSWCAP3 SWCAP3 VSS pwl 0.09us 0V 0.1us {AVDD} 

* VSWDRAIN1 SWDRAIN1 VSS dc {AVDD}
* VSWDRAIN2 SWDRAIN2 VSS dc {AVDD}
* VSWDRAIN2 SWDRAIN3 VSS dc {AVDD}
VSWDRAIN1 SWDRN1 VSS dc 0
VSWDRAIN2 SWDRN2 VSS dc 0
VSWDRAIN3 SWDRN3 VSS dc 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .option savecurrents
* .save all

* .save v(iout)
* .save v(xdut.x1.pbias) v(xdut.x1.nbias)
* .save v(b0) v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) v(b7) 
* .save v(bt)
* .save v(xdut.x1.b0_n) v(xdut.x1.b1_n) v(xdut.x1.b2_n) v(xdut.x1.b3_n) v(xdut.x1.b4_n)
* .save v(xdut.x1.v0) v(xdut.x1.v1) v(xdut.x1.v2) v(xdut.x1.v3) v(xdut.x1.v4)
* .save v(xdut.x1.vctrl) v(xdut.x1.vctrl_b)
* .save v(vdd) v(vss) v(sleep)

.save 
+ v(b0) v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) v(b7) v(bt)
+ v(xdut.iout)
+ v(xdut.src1) v(xdut.src2) v(xdut.src3)
+ v(xdut.vref) v(vout)
+ v(v1) 
+ v(xdut.v1a) v(xdut.v1b) 
+ v(v2) 
+ v(xdut.v2a) v(xdut.v2b) v(xdut.v2c)
+ v(xdut.x1.ctl) v(xdut.x1.ctlb) v(xdut.x1.vt)
+ v(vss) v(vdd) v(slp)
+ i(v.xdut.v1)
+ clock_frequency
+ duty_cycle
* + v(xdut.r1) v(xdut.r2)
* + v(xdut.x1.b0_n) v(xdut.x1.b1_n) v(xdut.x1.b2_n) v(xdut.x1.b3_n) v(xdut.x1.b4_n) v(xdut.x1.b5_n) v(xdut.x1.b6_n) v(xdut.x1.b7_n) v(xdut.x1.bt_n)
* + v(xdut.x1.pbias) v(xdut.x1.nbias) 
* + v(xdut.x1.v0) v(xdut.x1.v1) v(xdut.x1.v2) v(xdut.x1.v3) v(xdut.x1.v4) v(xdut.x1.v5) v(xdut.x1.v6) v(xdut.x1.v7)
* + v(SWBRN1) v(SWBRN2) v(SWBRN3) v(SWBGR1) v(SWBGR2) v(SWCAP1) v(SWCAP2) v(SWCAP3) v(SWDRN1) v(SWDRN2) v(SWDRN3)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

option temp = $&circuit_temperature

optran 0 0 0 1ns 1us 0

set fend = .raw
set clk_freq = {$&clock_frequency}
set clk_per = {1/clk_freq}
set cir_temp = {$&circuit_temperature}
set dcycle = {$&duty_cycle}
set vsup = {$&voltage_supply}

tran 1ns $&simulation_length 1ps
write {cicname}_temperature{$cir_temp}celsius_frequency{$clk_freq}mhz_dutycycle{$dcycle}percent_vdd{$vsup}volt{$fend}
* write

echo Circuit temperature: $cir_temp Celsius.
echo Simulation lenght: $&simulation_length seconds.
echo Clock frequency of finetuning signal: {$clk_freq} Mega Hertz, and clock periode is: {$clk_per} micro seconds.
echo Duty cycle of fine tuning signal: {$dcycle} %.
echo Supply voltage (VDD): {$vsup} Volt.
echo Circuit process corners: {cicname}.

* foreach vtemp -40 0 27 125
* 	reset
* 	option temp=$vtemp
* 	op
* 	tran 1ns $simulation_length 1ps
* 	write {cicname}_$vtemp$fend
* end

quit

.endc

.end