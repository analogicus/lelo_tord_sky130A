*Automatic generated instance fron ../../tech/scripts/genxdut dig
adut [cmp
+ rst
+ ]
+ [rst_out
+ sel_cap1
+ sel_cap2
+ b.7
+ b.6
+ b.5
+ b.4
+ b.3
+ b.2
+ b.1
+ b.0
+ ] null dut
.model dut d_cosim simulation="../dig.so" delay=10p

* Inputs
Rsvi0 cmp 0 1G
Rsvi1 rst 0 1G

* Outputs
Rsvi2 rst_out 0 1G
Rsvi3 sel_cap1 0 1G
Rsvi4 sel_cap2 0 1G
Rsvi5 b.7 0 1G
Rsvi6 b.6 0 1G
Rsvi7 b.5 0 1G
Rsvi8 b.4 0 1G
Rsvi9 b.3 0 1G
Rsvi10 b.2 0 1G
Rsvi11 b.1 0 1G
Rsvi12 b.0 0 1G

.save v(rst_out)

.save v(sel_cap1)

.save v(sel_cap2)

E_STATE_b dec_b 0 value={( 0 
+ + 128*v(b.7)/AVDD
+ + 64*v(b.6)/AVDD
+ + 32*v(b.5)/AVDD
+ + 16*v(b.4)/AVDD
+ + 8*v(b.3)/AVDD
+ + 4*v(b.2)/AVDD
+ + 2*v(b.1)/AVDD
+ + 1*v(b.0)/AVDD
+)/1000}
.save v(dec_b)

