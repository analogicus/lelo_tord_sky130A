magic
tech sky130A
timestamp 1770505916
<< locali >>
rect 1934 5791 7016 5794
rect 1934 5701 2039 5791
rect 2129 5786 3839 5791
rect 2129 5701 2939 5786
rect 1934 5698 2939 5701
rect 1844 4844 1940 5698
rect 2420 4847 2516 5698
rect 1820 3994 1916 4483
rect 2420 3994 2516 4477
rect 2744 4044 2840 5698
rect 3029 5701 3839 5786
rect 3929 5786 5639 5791
rect 3929 5701 4739 5786
rect 3029 5698 4739 5701
rect 3320 4044 3416 5698
rect 3644 4044 3740 5698
rect 4220 4044 4316 5698
rect 4544 4044 4640 5698
rect 4829 5701 5639 5786
rect 5729 5786 7016 5791
rect 5729 5701 6539 5786
rect 4829 5698 6539 5701
rect 5120 4045 5216 5698
rect 5444 4044 5540 5698
rect 6020 4044 6116 5698
rect 6344 4844 6440 5698
rect 6629 5698 7016 5786
rect 6920 4844 7016 5698
rect 6344 3996 6440 4487
rect 6920 3996 7016 4482
rect 6344 3994 7016 3996
rect 1494 3993 7016 3994
rect 1494 3991 6539 3993
rect 1494 3901 2039 3991
rect 2129 3903 6539 3991
rect 6629 3903 7016 3993
rect 2129 3901 7016 3903
rect 1494 3900 7016 3901
rect 1494 3898 6441 3900
rect 1494 3535 6115 3898
rect -156 3505 6115 3535
rect -156 3205 2840 3505
rect -156 3204 1637 3205
rect -156 2696 -60 3204
rect 420 2696 640 3204
rect -156 2606 39 2696
rect 129 2606 640 2696
rect -156 2600 640 2606
rect 544 2296 640 2600
rect 544 2207 739 2296
rect 1120 2296 1340 3204
rect 1820 2296 2840 3205
rect 3320 2296 3740 3505
rect 4220 2296 4640 3505
rect 5120 2296 5540 3505
rect 6019 3484 6115 3505
rect 6019 3418 6116 3484
rect 6020 2296 6116 3418
rect 829 2292 6116 2296
rect 829 2207 1439 2292
rect 544 2202 1439 2207
rect 1529 2202 6116 2292
rect 544 2200 6116 2202
<< viali >>
rect 1844 5698 1934 5794
rect 2039 5701 2129 5791
rect 1260 5416 1380 5530
rect 2939 5696 3029 5786
rect 3839 5701 3929 5791
rect 4739 5696 4829 5786
rect 5639 5701 5729 5791
rect 6539 5696 6629 5786
rect 2039 3901 2129 3991
rect 6539 3903 6629 3993
rect 1260 3682 1374 3802
rect 39 2606 129 2696
rect 739 2207 829 2297
rect 1439 2202 1529 2292
<< metal1 >>
rect 1841 5794 1937 5800
rect 1259 5698 1844 5794
rect 1934 5698 1937 5794
rect 1260 5533 1380 5698
rect 1841 5692 1937 5698
rect 2036 5791 2132 5797
rect 2036 5701 2039 5791
rect 2129 5701 2132 5791
rect 1254 5530 1386 5533
rect 1254 5416 1260 5530
rect 1380 5416 1386 5530
rect 1254 5413 1386 5416
rect 1972 4923 2004 5638
rect 2036 5112 2132 5701
rect 2936 5786 3032 5792
rect 2936 5696 2939 5786
rect 3029 5696 3032 5786
rect 1972 4888 2004 4891
rect 1972 4282 2004 4285
rect 1972 4171 2004 4250
rect 2036 3991 2132 4408
rect 2228 4282 2324 5644
rect 2228 4250 2259 4282
rect 2291 4250 2324 4282
rect 2228 4084 2324 4250
rect 2872 4923 2904 5607
rect 2872 4115 2904 4891
rect 2936 4312 3032 5696
rect 3836 5791 3932 5797
rect 3836 5701 3839 5791
rect 3929 5701 3932 5791
rect 3128 4923 3224 5639
rect 3128 4891 3158 4923
rect 3190 4891 3224 4923
rect 2036 3901 2039 3991
rect 2129 3901 2132 3991
rect 2036 3895 2132 3901
rect 1257 3802 1377 3808
rect 636 3682 1260 3802
rect 1374 3682 1377 3802
rect 636 3460 756 3682
rect 1257 3676 1377 3682
rect 3128 3701 3224 4891
rect 3772 4840 3804 5602
rect 3772 4120 3804 4808
rect 3836 4312 3932 5701
rect 4736 5786 4832 5792
rect 4736 5696 4739 5786
rect 4829 5696 4832 5786
rect 4028 4923 4124 5639
rect 4028 4891 4056 4923
rect 4088 4891 4124 4923
rect 4028 3701 4124 4891
rect 4672 4923 4704 5587
rect 4672 4084 4704 4891
rect 4736 4312 4832 5696
rect 5636 5791 5732 5797
rect 5636 5701 5639 5791
rect 5729 5701 5732 5791
rect 4928 4840 5024 5639
rect 4928 4808 4959 4840
rect 4991 4808 5024 4840
rect 3128 3605 4124 3701
rect -28 3443 1403 3460
rect -28 3340 1404 3443
rect -28 2784 4 3340
rect 36 2696 132 3108
rect 228 2784 324 3340
rect 36 2606 39 2696
rect 129 2606 132 2696
rect 36 2600 132 2606
rect 672 2484 704 3340
rect 736 2297 832 3108
rect 736 2207 739 2297
rect 829 2207 832 2297
rect 736 2201 832 2207
rect 928 2166 1024 2852
rect 1372 2384 1404 3340
rect 1436 2292 1532 3108
rect 2872 2925 2904 3443
rect 2869 2893 2872 2925
rect 2904 2893 2907 2925
rect 1436 2202 1439 2292
rect 1529 2202 1532 2292
rect 1436 2196 1532 2202
rect 1628 2166 1724 2848
rect 2872 2384 2904 2893
rect 2936 2166 3032 3408
rect 3128 2384 3224 3605
rect 3772 2925 3804 3443
rect 3772 2384 3804 2893
rect 3836 2166 3932 3408
rect 4028 2384 4124 3605
rect 4928 3699 5024 4808
rect 5572 4840 5604 5592
rect 5572 4120 5604 4808
rect 5636 4312 5732 5701
rect 6536 5786 6632 5792
rect 6536 5696 6539 5786
rect 6629 5696 6632 5786
rect 5828 4840 5924 5644
rect 6472 4844 6504 5571
rect 6536 5112 6632 5696
rect 5828 4808 5859 4840
rect 5891 4808 5924 4840
rect 5828 3699 5924 4808
rect 6469 4840 6509 4844
rect 6469 4808 6472 4840
rect 6504 4808 6509 4840
rect 6469 4804 6509 4808
rect 6471 4282 6503 4285
rect 6471 4247 6503 4250
rect 6536 3993 6632 4408
rect 6728 4084 6824 5649
rect 6536 3903 6539 3993
rect 6629 3903 6632 3993
rect 6536 3897 6632 3903
rect 4928 3603 5924 3699
rect 4672 2915 4704 3438
rect 4669 2883 4672 2915
rect 4704 2883 4707 2915
rect 4672 2384 4704 2883
rect 4736 2166 4832 3408
rect 4928 2384 5024 3603
rect 5572 2915 5604 3435
rect 5572 2384 5604 2883
rect 5636 2166 5732 3408
rect 5828 2384 5924 3603
rect 928 2070 5732 2166
<< via1 >>
rect 1972 4891 2004 4923
rect 1972 4250 2004 4282
rect 2259 4250 2291 4282
rect 2872 4891 2904 4923
rect 3158 4891 3190 4923
rect 3772 4808 3804 4840
rect 4056 4891 4088 4923
rect 4672 4891 4704 4923
rect 4959 4808 4991 4840
rect 2872 2893 2904 2925
rect 3772 2893 3804 2925
rect 5572 4808 5604 4840
rect 5859 4808 5891 4840
rect 6472 4808 6504 4840
rect 6471 4250 6503 4282
rect 4672 2883 4704 2915
rect 5572 2883 5604 2915
<< metal2 >>
rect 1969 4891 1972 4923
rect 2004 4891 2872 4923
rect 2904 4891 3158 4923
rect 3190 4891 4056 4923
rect 4088 4891 4672 4923
rect 4704 4891 4707 4923
rect 6469 4840 6509 4844
rect 3769 4808 3772 4840
rect 3804 4808 4959 4840
rect 4991 4808 5572 4840
rect 5604 4808 5859 4840
rect 5891 4808 6472 4840
rect 6504 4808 6509 4840
rect 6469 4804 6509 4808
rect 1969 4250 1972 4282
rect 2004 4250 2259 4282
rect 2291 4250 6471 4282
rect 6503 4250 6506 4282
rect 2872 2925 2904 2928
rect 2904 2893 3772 2925
rect 3804 2893 3807 2925
rect 4672 2915 4704 2918
rect 5559 2915 5611 2923
rect 2872 2890 2904 2893
rect 4704 2883 5572 2915
rect 5604 2883 5611 2915
rect 4672 2880 4704 2883
rect 5559 2877 5611 2883
use JNWATR_NCH_4C5F0  xa8<0> ~/pro/aicex/ip/lelo_tord_sky130A/design/JNW_ATR_SKY130A
timestamp 1770500839
transform 1 0 2792 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa8<1>
timestamp 1770500839
transform 1 0 2792 0 1 3064
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa8<2>
timestamp 1770500839
transform 1 0 3692 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa8<3>
timestamp 1770500839
transform 1 0 3692 0 1 3064
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa9<0>
timestamp 1770500839
transform 1 0 5492 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa9<1>
timestamp 1770500839
transform 1 0 5492 0 1 3064
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa9<2>
timestamp 1770500839
transform 1 0 4592 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xa9<3>
timestamp 1770500839
transform 1 0 4592 0 1 3064
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb12
timestamp 1770500839
transform 1 0 -108 0 1 2764
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb13<0>
timestamp 1770500839
transform 1 0 592 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb13<1>
timestamp 1770500839
transform 1 0 592 0 1 2764
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb13<2>
timestamp 1770500839
transform 1 0 1292 0 1 2364
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb13<3>
timestamp 1770500839
transform 1 0 1292 0 1 2764
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xc10
timestamp 1770500839
transform 1 0 1892 0 1 4064
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xc11
timestamp 1770500839
transform 1 0 6392 0 1 4064
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd2<0> ~/pro/aicex/ip/lelo_tord_sky130A/design/LELO_TORD_SKY130A/../JNW_ATR_SKY130A
timestamp 1770384003
transform 1 0 1892 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd2<1>
timestamp 1770384003
transform 1 0 1892 0 1 5264
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd3<0>
timestamp 1770384003
transform 1 0 2792 0 1 4064
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd3<1>
timestamp 1770384003
transform 1 0 2792 0 1 4464
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd3<2>
timestamp 1770384003
transform 1 0 2792 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd3<3>
timestamp 1770384003
transform 1 0 2792 0 1 5264
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd4<0>
timestamp 1770384003
transform 1 0 3692 0 1 4064
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd4<1>
timestamp 1770384003
transform 1 0 3692 0 1 4464
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd4<2>
timestamp 1770384003
transform 1 0 3692 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd4<3>
timestamp 1770384003
transform 1 0 3692 0 1 5264
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd5<0>
timestamp 1770384003
transform 1 0 4592 0 1 4064
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd5<1>
timestamp 1770384003
transform 1 0 4592 0 1 4464
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd5<2>
timestamp 1770384003
transform 1 0 4592 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd5<3>
timestamp 1770384003
transform 1 0 4592 0 1 5264
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd6<0>
timestamp 1770384003
transform 1 0 5492 0 1 4064
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd6<1>
timestamp 1770384003
transform 1 0 5492 0 1 4464
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd6<2>
timestamp 1770384003
transform 1 0 5492 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd6<3>
timestamp 1770384003
transform 1 0 5492 0 1 5264
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd7<0>
timestamp 1770384003
transform 1 0 6392 0 1 4864
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xd7<1>
timestamp 1770384003
transform 1 0 6392 0 1 5264
box -92 -64 668 464
use JNWTR_RPPO16  xr1 ~/pro/aicex/ip/lelo_tord_sky130A/design/LELO_TORD_SKY130A/../JNW_TR_SKY130A
timestamp 1770374940
transform 0 1 -200 -1 0 5736
box 0 0 2236 1720
<< labels >>
flabel metal1 s 2036 5164 2132 5204 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal1 s 2228 4084 2324 4124 0 FreeSans 200 0 0 0 VOUT_N
port 5 nsew signal bidirectional
flabel metal1 s 5572 2544 5604 2584 0 FreeSans 200 0 0 0 VIN
port 3 nsew signal bidirectional
flabel metal1 s 2872 2544 2904 2584 0 FreeSans 200 0 0 0 VIP
port 4 nsew signal bidirectional
flabel locali s 2744 2544 2840 2584 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional
flabel metal1 s 6728 4084 6824 4124 0 FreeSans 200 0 0 0 VOUT
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX -48 0 5900 8000
<< end >>
