*Automatic generated instance fron ../../tech/scripts/genxdut dac_v2
adut [clk
+ rst
+ ]
+ [b.3
+ b.2
+ b.1
+ b.0
+ count.2
+ count.1
+ count.0
+ ] null dut
.model dut d_cosim simulation="../dac_v2.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 rst 0 1G

* Outputs
Rsvi2 b.3 0 1G
Rsvi3 b.2 0 1G
Rsvi4 b.1 0 1G
Rsvi5 b.0 0 1G
Rsvi6 count.2 0 1G
Rsvi7 count.1 0 1G
Rsvi8 count.0 0 1G

E_STATE_b dec_b 0 value={( 0 
+ + 8*v(b.3)/AVDD
+ + 4*v(b.2)/AVDD
+ + 2*v(b.1)/AVDD
+ + 1*v(b.0)/AVDD
+)/1000}
.save v(dec_b)

E_STATE_count dec_count 0 value={( 0 
+ + 4*v(count.2)/AVDD
+ + 2*v(count.1)/AVDD
+ + 1*v(count.0)/AVDD
+)/1000}
.save v(dec_count)

