*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_dac_and_bgr.spi
#else
.include ../../../work/xsch/TB_dac_and_bgr.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10ps
.param AVDD = {vdda}

.param f_CLK = 2MegHz
.param T_CLK = {1/f_CLK}

.param TD = {T_CLK}
.param TR = {T_CLK/100}
.param TF = {TR}
.param PW = {T_CLK}
.param PER = {T_CLK}

* Time averaging duty cycle is given in percent (%)
.param dutycycle = 35
.param ratio = {dutycycle/100}

* Stepping Current out of DAC
.param step_start = 0.5us
.param step_length = 2.0us

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS   VSS   0    dc 0V
VDD   VDD   VSS  dc {AVDD}
VSLP  SLP VSS pwl 0.02us {AVDD} 0.03us 0V

* VB0  B0   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*8/16} {PER})
* VB1  B1   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*9/16} {PER})
* VB2  B2   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*10/16} {PER})
* VB3  B3   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*11/16} {PER})
* VB4  B4   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*12/16} {PER})
* VB5  B5   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*13/16} {PER})
* VB6  B6   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*14/16} {PER})
* VB7  B7   VSS  PULSE({AVDD} 0V {TD} {TR} {TF} {PW*15/16} {PER})

VB0  B0   VSS  dc pwl {step_start + 0*step_length} 0V {step_start + 0*step_length + 0.01us} {AVDD}
VB1  B1   VSS  dc pwl {step_start + 1*step_length} 0V {step_start + 1*step_length + 0.01us} {AVDD}
VB2  B2   VSS  dc pwl {step_start + 2*step_length} 0V {step_start + 2*step_length + 0.01us} {AVDD}
VB3  B3   VSS  dc pwl {step_start + 3*step_length} 0V {step_start + 3*step_length + 0.01us} {AVDD}
VB4  B4   VSS  dc pwl {step_start + 4*step_length} 0V {step_start + 4*step_length + 0.01us} {AVDD}
VB5  B5   VSS  dc pwl {step_start + 5*step_length} 0V {step_start + 5*step_length + 0.01us} {AVDD}
VB6  B6   VSS  dc pwl {step_start + 6*step_length} 0V {step_start + 6*step_length + 0.01us} {AVDD}
VB7  B7   VSS  dc pwl {step_start + 7*step_length} 0V {step_start + 7*step_length + 0.01us} {AVDD}

* VBT  BT   VSS  PULSE({AVDD} 0V {2*TD} {TR} {TF} {PW*ratio} {PER})
VBT  BT   VSS  PULSE(0V {AVDD} {2*TD} {TR} {TF} {PW*ratio} {PER})
* VBT  BT   VSS  DC 0V

VSWBRANCH1 SWBRN1 VSS dc {AVDD}
VSWBRANCH2 SWBRN2 VSS dc {AVDD}
VSWBRANCH3 SWBRN3 VSS dc {AVDD}
* VSWBRANCH1 SWBRN1 VSS dc 0
* VSWBRANCH2 SWBRN2 VSS dc 0
* VSWBRANCH3 SWBRN3 VSS dc 0

VSWBGR1 SWBGR1 VSS dc {AVDD}
VSWBGR2 SWBGR2 VSS dc {AVDD}
* VSWBGR1 SWBGR1 VSS dc 0
* VSWBGR2 SWBGR2 VSS dc 0

* VSWCAP1 SWCAP1 VSS dc {AVDD}
* VSWCAP2 SWCAP2 VSS dc {AVDD}
* VSWCAP3 SWCAP3 VSS dc {AVDD}
* VSWCAP1 SWCAP1 VSS dc 0
* VSWCAP2 SWCAP2 VSS dc 0
* VSWCAP3 SWCAP3 VSS dc 0
VSWCAP1 SWCAP1 VSS pwl 0.09us 0V 0.1us {AVDD} 
VSWCAP2 SWCAP2 VSS pwl 0.09us 0V 0.1us {AVDD} 
VSWCAP3 SWCAP3 VSS pwl 0.09us 0V 0.1us {AVDD} 

* VSWDRAIN1 SWDRAIN1 VSS dc {AVDD}
* VSWDRAIN2 SWDRAIN2 VSS dc {AVDD}
* VSWDRAIN2 SWDRAIN3 VSS dc {AVDD}
VSWDRAIN1 SWDRN1 VSS dc 0
VSWDRAIN2 SWDRN2 VSS dc 0
VSWDRAIN3 SWDRN3 VSS dc 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .option savecurrents
* .save all

* .save v(iout)
* .save v(xdut.x1.pbias) v(xdut.x1.nbias)
* .save v(b0) v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) v(b7) 
* .save v(bt)
* .save v(xdut.x1.b0_n) v(xdut.x1.b1_n) v(xdut.x1.b2_n) v(xdut.x1.b3_n) v(xdut.x1.b4_n)
* .save v(xdut.x1.v0) v(xdut.x1.v1) v(xdut.x1.v2) v(xdut.x1.v3) v(xdut.x1.v4)
* .save v(xdut.x1.vctrl) v(xdut.x1.vctrl_b)
* .save v(vdd) v(vss) v(sleep)

.save 
+ v(b0) v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) v(b7) v(bt)
+ v(SWBRN1) v(SWBRN2) v(SWBRN3) v(SWBGR1) v(SWBGR2) v(SWCAP1) v(SWCAP2) v(SWCAP3) v(SWDRN1) v(SWDRN2) v(SWDRN3)
+ v(xdut.iout)
+ v(xdut.src1) v(xdut.src2) v(xdut.src3)
+ v(xdut.vref) v(vout)
+ v(v1) 
+ v(xdut.v1a) v(xdut.v1b) 
+ v(v2) 
+ v(xdut.v2a) v(xdut.v2b) v(xdut.v2c)
+ v(xdut.r1) v(xdut.r2)
+ v(xdut.x1.ctl) v(xdut.x1.ctlb) v(xdut.x1.vt)
+ v(xdut.x1.b0_n) v(xdut.x1.b1_n) v(xdut.x1.b2_n) v(xdut.x1.b3_n) v(xdut.x1.b4_n) v(xdut.x1.b5_n) v(xdut.x1.b6_n) v(xdut.x1.b7_n) v(xdut.x1.bt_n)
+ v(xdut.x1.v0) v(xdut.x1.v1) v(xdut.x1.v2) v(xdut.x1.v3) v(xdut.x1.v4) v(xdut.x1.v5) v(xdut.x1.v6) v(xdut.x1.v7)
+ v(xdut.x1.pbias) v(xdut.x1.nbias) 
+ v(vss) v(vdd) v(slp)
+ i(v.xdut.v1)

*test

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1ns 1us 0


set simulation_length = 16.5us

tran 1ns $simulation_length 1ps
write

set fend = .raw
foreach vtemp -45 -25 0 25 50 75 100 125
	option temp=$vtemp
	tran 1ns $simulation_length 1ps
	write {cicname}_$vtemp$fend
end

quit


.endc

.end