*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_dig_ctrl_lpe.spi
#else
.include ../../../work/xsch/TB_dig_ctrl.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

* Analog supply voltage given in Volts (V)
.param AVDD = {vdda}
.csparam voltage_supply_csparam = {vdda}

* Circuit temperature given in degrees Celsius (C)
.param circuit_temperature = 27
.csparam circuit_temperature_csparam = {circuit_temperature}

* Time averaging finetuning duty cycle is given in percent (%)
.param finetuning_dutycycle = 40
.csparam finetuning_dutycycle_csparam = {finetuning_dutycycle}

.param ratio = finetuning_dutycycle/100

* finetuning_frequency = 2 MHz => finetuning_periode = 0.5 us
* finetuning_frequency = 1 MHz => finetuning_periode = 1.0 us
.param finetuning_frequency = 1
.csparam finetuning_frequency_csparam = {finetuning_frequency}

.param finetuning_frequency_MHz = finetuning_frequency*1MegHz
.param finetuning_periode = 1/finetuning_frequency_MHz
.param TD = finetuning_periode
.param TR = finetuning_periode/100
.param TF = TR
.param PW = finetuning_periode
.param PER = finetuning_periode

* Stepping Current out of DAC
.param step_start = 25us
.param step_length = 5.0us

* .csparam simulation_length_csparam = {step_start + 16*step_length}
.csparam simulation_length_csparam = {step_start + 7*step_length}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0    dc  0V
VDD  VDD  VSS  dc  {AVDD}
VSLP SLP  VSS  pwl 0.02us {AVDD} 0.03us 0V

VCLK CLK  VSS  PULSE(0V {AVDD} {2*TD} {TR} {TF} {PW*ratio} {PER})
VRST RESET VSS PWL 30us 0V 31us {AVDD} 39us {AVDD} 40us 0V

* VB1  B1   VSS  dc pwl {step_start + 1*step_length}  0V {step_start + 1*step_length  + 0.01us} {AVDD}
* VB2  B2   VSS  dc pwl {step_start + 2*step_length}  0V {step_start + 2*step_length  + 0.01us} {AVDD}
* VB3  B3   VSS  dc pwl {step_start + 3*step_length}  0V {step_start + 3*step_length  + 0.01us} {AVDD}
VB4  B4   VSS  dc pwl {step_start + 4*step_length}  0V {step_start + 4*step_length  + 0.01us} {AVDD}
VB5  B5   VSS  dc pwl {step_start + 5*step_length}  0V {step_start + 5*step_length  + 0.01us} {AVDD}
VB6  B6   VSS  dc pwl {step_start + 6*step_length}  0V {step_start + 6*step_length  + 0.01us} {AVDD}
* VB7  B7   VSS  dc pwl {step_start + 7*step_length}  0V {step_start + 7*step_length  + 0.01us} {AVDD}
* VB8  B8   VSS  dc pwl {step_start + 8*step_length}  0V {step_start + 8*step_length  + 0.01us} {AVDD}
* VB9  B9   VSS  dc pwl {step_start + 9*step_length}  0V {step_start + 9*step_length  + 0.01us} {AVDD}
* VB10 B10  VSS  dc pwl {step_start + 10*step_length} 0V {step_start + 10*step_length + 0.01us} {AVDD}
* VB11 B11  VSS  dc pwl {step_start + 11*step_length} 0V {step_start + 11*step_length + 0.01us} {AVDD}
* VB12 B12  VSS  dc pwl {step_start + 12*step_length} 0V {step_start + 12*step_length + 0.01us} {AVDD}
* VB13 B13  VSS  dc pwl {step_start + 13*step_length} 0V {step_start + 13*step_length + 0.01us} {AVDD}
* VB14 B14  VSS  dc pwl {step_start + 14*step_length} 0V {step_start + 14*step_length + 0.01us} {AVDD}
* VB15 B15  VSS  dc pwl {step_start + 15*step_length} 0V {step_start + 15*step_length + 0.01us} {AVDD}

VB1  B1   VSS  dc {AVDD}
VB2  B2   VSS  dc {AVDD}
VB3  B3   VSS  dc {AVDD}
* VB4  B4   VSS  dc {AVDD}
* VB5  B5   VSS  dc {AVDD}
* VB6  B6   VSS  dc 0V
VB7  B7   VSS  dc 0V
VB8  B8   VSS  dc 0V
VB9  B9   VSS  dc 0V
VB10  B10   VSS  dc 0V
VB11  B11   VSS  dc 0V
VB12  B12   VSS  dc 0V
VB13  B13   VSS  dc 0V
VB14  B14   VSS  dc 0V
VB15  B15   VSS  dc 0V

VBT  BT   VSS  PULSE(0V {AVDD} {2*TD} {TR} {TF} {PW*ratio} {PER})

VSWBRANCH1 SWBRN1 VSS dc {AVDD}
VSWBRANCH2 SWBRN2 VSS dc {AVDD}
VSWBRANCH3 SWBRN3 VSS dc {AVDD}

VSWBGR1 SWBGR1 VSS dc 0V
VSWBGR2 SWBGR2 VSS dc 0V

VSWCAP1 SWCAP1 VSS dc {AVDD}
VSWCAP2 SWCAP2 VSS dc {AVDD}
VSWCAP3 SWCAP3 VSS dc {AVDD}

VSWDRAIN1 SWDRN1 VSS dc 0V
VSWDRAIN2 SWDRN2 VSS dc 0V
VSWDRAIN3 SWDRN3 VSS dc 0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names (Do not use the letter t or any number to replace x in VBx, as they have already most likely been used)
VBa b.0 b<0> dc 0
VBb b.1 b<1> dc 0
VBc b.2 b<2> dc 0
VBd b.3 b<3> dc 0
VBe b.4 b<4> dc 0

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .save all

.save 
+ v(b1) v(b2) v(b3)  v(b4)  v(b5)  v(b6)  v(b7)
+ v(b8) v(b9) v(b10) v(b11) v(b12) v(b13) v(b14) v(b15) 
+ v(bt)
+ v(xdut.iout)
+ v(xdut.src1) v(xdut.src2) v(xdut.src3)
+ v(xdut.vref) v(vout)
+ v(cmp)
+ v(v1) 
+ v(xdut.v1a) v(xdut.v1b) 
+ v(v2) 
+ v(xdut.v2a) v(xdut.v2b) v(xdut.v2c)
+ v(xdut.x1.ctl) v(xdut.x1.ctlb) v(xdut.x1.vt)
+ v(vss) v(vdd) v(slp)
+ i(v.xdut.v1)
+ i(vss) i(vdd)
* + v(xdut.r1) v(xdut.r2)
* + v(xdut.x1.b1_n) v(xdut.x1.b2_n) v(xdut.x1.b3_n)  v(xdut.x1.b4_n)  v(xdut.x1.b5_n)  v(xdut.x1.b6_n)  v(xdut.x1.b7_n)
* + v(xdut.x1.b8_n) v(xdut.x1.b9_n) v(xdut.x1.b10_n) v(xdut.x1.b11_n) v(xdut.x1.b12_n) v(xdut.x1.b13_n) v(xdut.x1.b14_n) v(xdut.x1.b15_n)
* + v(xdut.x1.bt_n)
* + v(xdut.x1.pbias) v(xdut.x1.nbias) 
* + v(xdut.x1.v0) v(xdut.x1.v1) v(xdut.x1.v2) v(xdut.x1.v3) v(xdut.x1.v4) v(xdut.x1.v5) v(xdut.x1.v6) v(xdut.x1.v7)
* + v(SWBRN1) v(SWBRN2) v(SWBRN3) v(SWBGR1) v(SWBGR2) v(SWCAP1) v(SWCAP2) v(SWCAP3) v(SWDRN1) v(SWDRN2) v(SWDRN3)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

set vsupply = {$&voltage_supply_csparam}
set cirtemp = {$&circuit_temperature_csparam}
set clkfreq = {$&finetuning_frequency_csparam}
set clkper = {1/$clkfreq}
set dcycle = {$&finetuning_dutycycle_csparam}
set simlen = {$&simulation_length_csparam}

echo $vsupply
echo $cirtemp
echo $clkfreq
echo $clkper
echo $dcycle
echo $simlen

* temperature options: -40 -20 0 27 60 90 125
* dutycycle options:  10 20 30 40 50 60 70 80 90

set fend = .raw
foreach cirtemp 27
	foreach clkfreq 1
		foreach dcycle 50
			option temp = $cirtemp
			alterparam finetuning_frequency = {$clkfreq}
			alterparam finetuning_dutycycle = {$dcycle}
            reset

			* if your netlist uses derived params like ratio from dutycycle,
			* they will re-evaluate automatically as long as they are expressions:
			*   .param clkper = {1/clkfreq}
			*   .param ratio = {dcycle/100}

			let clkper = {1/$clkfreq}

			echo ------------------------------------------------------------
			echo VDD: $vsupply V
			echo Temperature: $cirtemp C
			echo Finetuning frequency: $clkfreq MHz, Period: $clkper us
			echo Duty cycle: $dcycle %
			echo Corner: {cicname}
			echo Simulation lenght: $simlen seconds.
			echo ------------------------------------------------------------

			optran 0 0 0 1ns 1us 0
			tran 1ns $simlen 1ps

			write {cicname}_temperature{$cirtemp}celsius_frequency{$clkfreq}mhz_dutycycle{$dcycle}percent_vdd{$vsupply}volt{$fend}

			*
			* This last part used to be in tran.meas, but was moved to ensure all simulations are written to .out-files
			*

			load {cicname}_temperature{$cirtemp}celsius_frequency{$clkfreq}mhz_dutycycle{$dcycle}percent_vdd{$vsupply}volt{$fend}

			let v(x1.vt) = v(xdut.x1.vt)
			let v(x1.ctl) = v(xdut.x1.ctl)
			let v(x1.ctlb) = v(xdut.x1.ctlb)

			let v(iout) = v(xdut.iout)

			let v(src1) = v(xdut.src1) 
			let v(src2) = v(xdut.src2)
			let v(src3) = v(xdut.src3)
			let v(v1a) = v(xdut.v1a)
			let v(v1b) = v(xdut.v1b)
			let v(v2a) = v(xdut.v2a)
			let v(v2b) = v(xdut.v2b)
			let v(v2c) = v(xdut.v2c)
			let v(vref) = v(xdut.vref)

			set fend = .out
			set wr_singlescale
			set wr_vecnames
			option numdgt = 5
			echo writing to {cicname}_temperature{$cirtemp}celsius_frequency{$clkfreq}mhz_dutycycle{$dcycle}percent_vdd{$vsupply}volt{$fend}
			wrdata {cicname}_temperature{$cirtemp}celsius_frequency{$clkfreq}mhz_dutycycle{$dcycle}percent_vdd{$vsupply}volt{$fend}
            + v(b1) v(b2) v(b3) v(b4) v(b5) v(b6) v(b7) 
            + v(b8) v(b9) v(b10) v(b11) v(b12) v(b13) v(b14) v(b15) 
            + v(bt)
			+ v(iout)
			+ v(src1) v(src2) v(src3)
			+ v(vref) v(vout)
            + v(cmp)
			+ v(v1)
			+ v(v1a) v(v1b) 
			+ v(v2) 
			+ v(v2a) v(v2b) v(v2c)
			+ v(x1.ctl) v(x1.ctlb) v(x1.vt)
			+ v(vss) v(vdd) v(slp)
			+ i(v.xdut.v1)
			+ i(vdd) i(vss)
			+ v(dec_b)
		end
	end
end

quit

.endc

.end
