*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_inverters_lpe.spi
#else
.include ../../../work/xsch/TB_inverters.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0   dc  0
VDD VDD VSS dc  {AVDD}
V1  in1 vss pwl 0ns 0V 20ns {AVDD}
V2  in2 vss pwl 0ns 0V 20ns {AVDD}
V3  in3 vss pwl 0ns 0V 20ns {AVDD}
V4  in4 vss pwl 0ns 0V 20ns {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .option savecurrents
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1ns 1us 0


tran 1ns 20ns 1ps
write
quit


.endc

.end
