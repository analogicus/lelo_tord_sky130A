*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/cmp_v2_lpe.spi
#else
.include ../../../work/xsch/cmp_v2.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0    dc 0
VDD  VDD  VSS  dc {AVDD}
*VIP  VIP  VSS  pwl 0s 0V 0.1us 0V 1us {AVDD} 1.1us 0V 2us {AVDD} 2.1us 0V 3us {AVDD} 3.1us 0V
*VIN  VIN  VSS  dc 0.9V
VIP  VIP  VSS  pwl 0s 0V 1us {AVDD} 2us 0V 3us {AVDD} 4us 0V 4.5us {AVDD}
VIN  VIN  VSS  pwl 0s {AVDD} 1us 0V 2us {AVDD} 3us 0V 4us {AVDD} 4.5us 0V
*Vip  vip   VSS   pwl 0 0.89 1u 0.91 2u 0.89 3u 0.91 4u 0.89
*Vin  vin   VSS   pwl 0 0.91 1u 0.89 2u 0.91 3u 0.89 4u 0.91
*VIP VIP VSS SIN(0.9V 0.9V 1MEG 0s 0)
*VIN VIN VSS SIN(0.9V 0.9V 1MEG 0.5us 0)

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 5u 1p
write
quit


.endc

.end
