*Automatic generated instance fron ../../tech/scripts/genxdut digtotime
adut [clk
+ rst
+ ]
+ [d.3
+ d.2
+ d.1
+ d.0
+ count.2
+ count.1
+ count.0
+ ] null dut
.model dut d_cosim simulation="../digtotime.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 rst 0 1G

* Outputs
Rsvi2 d.3 0 1G
Rsvi3 d.2 0 1G
Rsvi4 d.1 0 1G
Rsvi5 d.0 0 1G
Rsvi6 count.2 0 1G
Rsvi7 count.1 0 1G
Rsvi8 count.0 0 1G

E_STATE_d dec_d 0 value={( 0 
+ + 8*v(d.3)/AVDD
+ + 4*v(d.2)/AVDD
+ + 2*v(d.1)/AVDD
+ + 1*v(d.0)/AVDD
+)/1000}
.save v(dec_d)

E_STATE_count dec_count 0 value={( 0 
+ + 4*v(count.2)/AVDD
+ + 2*v(count.1)/AVDD
+ + 1*v(count.0)/AVDD
+)/1000}
.save v(dec_count)

