*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bias_lpe.spi
#else
.include ../../../work/xsch/bias.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param delay = 10ns
.param rise = 1ns
.param width = 100ns
.param fall = 1ns

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0   dc 0
VDD VDD VSS dc {AVDD}
VSLEEP SLEEP VSS pwl {delay} 0V {delay+rise} {AVDD} {delay+rise+width} {AVDD} {delay+rise+width+fall} 0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents

*.save v(xdut.v1) v(xdut.v2) v(xdut.v3) v(xdut.v4) v(xdut.v5) v(xdut.v6)
*.save v(pbias)
*.save v(nbias)
*.save v(sleep)
*.save v(vdd) v(vss)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1ns 1us 0


tran 1ns 200ns 1ps
write
quit


.endc

.end
