*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bias_1p2u_lpe.spi
#else
.include ../../../work/xsch/bias_1p2u.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

.param delay = 10ns
.param rise = 1ns
.param width = 100ns
.param fall = 1ns

.param simulation_length = 400ns
* .param simulation_length = {delay + rise + width + fall + 200ns}

.csparam sim_len_csparam = {simulation_length}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0   dc 0V
VDD VDD VSS dc {AVDD}
* VSLEEP SLEEP VSS pwl {delay} 0V {delay+rise} {AVDD} {delay+rise+width} {AVDD} {delay+rise+width+fall} 0V
VSLEEP SLEEP VSS dc 0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

set sim_length = {$&sim_len_csparam}
echo $sim_length

optran 0 0 0 1ns 1us 0


tran 1ns $sim_length 1ps
write
quit


.endc

.end
