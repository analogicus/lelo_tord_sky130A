*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_tmp_core_and_cmp_lpe.spi
#else
.include ../../../work/xsch/TB_tmp_core_and_cmp.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD     VDD    VSS dc {AVDD}
IPTAT   VSS    IPTAT dc 750nA
*VSEL_C1 SEL_C1 VSS pulse(0V {AVDD} 1us 1ns 1ns 430ns 860ns)
*VSEL_C2 SEL_C2 VSS pulse({AVDD} 0V 1us 1ns 1ns 430ns 860ns)
*VRST    RST    VSS pwl 0s {AVDD} 0.9us {AVDD} 1us 0V 9us 0V 9.1us {AVDD} 9.2us {VDDA} 9.3us 0V
*VRST    RST    VSS pulse({AVDD} 0V 1us 10ns 10ns 1.9us 2us)
VRST    RST    VSS pwl 0.9us {AVDD} 1us 0V 8.5us 0V 8.6us {AVDD} 9.4us {AVDD} 9.5us 0V
VSS     VSS    0   dc 0V
VREF    REF    VSS dc 1.0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names
VB1 b.1 b<1> dc 0
VB2 b.2 b<2> dc 0
VB3 b.3 b<3> dc 0
VB4 b.4 b<4> dc 0
VB5 b.5 b<5> dc 0
VB6 b.6 b<6> dc 0
VB7 b.7 b<7> dc 0

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.option savecurrents
*.save all

* Save the voltages 
.save v(VDD)
.save v(VSS)
.save v(IPTAT)
*.save v(SEL_C1)
*.save v(SEL_C2)
.save v(RST)
.save v(REF)
.save v(CMP)
.save v(xdut.vptat)
.save v(xdut.x1.vcap1)
.save v(xdut.x1.vcap2)

.save v(b.7) v(b.6) v(b.5) v(b.4) v(b.3) v(b.2) v(b.1) v(b.0)

* Save the currents
*.save i(VDD)
*.save i(VSS)
*.save i(IPTAT)
*.save i(VSEL_C1)
*.save i(VSEL_C2)
*.save i(VRST)
*.save i(VREF)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

* Initial conditions (IC)
*ic v(iptat)=0 v(rst)=0

optran 0 0 0 1ns 10us 0


tran 1ns 30us
write
quit


.endc

.end
