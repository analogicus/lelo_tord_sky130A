*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_TORD_lpe.spi
.csparam schematic_or_layout = 8
#else
.include ../../../work/xsch/LELO_TORD.spice
.csparam schematic_or_layout = 9
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param CM = {AVDD/2} 

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0   DC 0V
VDD VDD VSS DC {AVDD}

VIP VIP VSS DC 0.9V AC 1V SIN(0.9V 10uV 100kHz)
VIN VIN VSS DC 0.9V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


echo begining transient analysis simulation

optran 0 0 0 1ns 10us 0
tran 1ns 10us 1ps
write {cicname}.raw


* Force ASCII format for raw file (human readable)
set filetype=ascii
let sch_or_lay = {$&schematic_or_layout}
write circuit_view.raw sch_or_lay

reset

* Reset to binary for efficiency
set filetype=binary


echo beginning ac analysis simulation

op
ac dec 100 1Hz 100MegHz
write {cicname}_ac.raw


* echo beginning dc analysis simulation

* dc vip 0.9V 1.1V 1mV
* write {cicname}_dc.raw

quit

.endc

.end

