*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/cmp_lpe.spi
#else
.include ../../../work/xsch/cmp.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param CM = {AVDD/2} 

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0   DC 0V
VDD VDD VSS DC {AVDD}

VIP VIP VSS DC 0.9V AC 1V SIN(0.9V 100uV 100kHz)
VIN VIN VSS DC 0.9V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1ns 10us 0

echo beginning tranisent analysis simulation

tran 1ns 11us 1ps
write {cicname}.raw

echo beginning ac analysis simulation

ac dec 100 1Hz 1GHz
write {cicname}_ac.raw

* echo beginning dc analysis simulation

* dc vip 0.9V 1.1V 1mV
* write {cicname}_dc.raw

quit

.endc

.end

