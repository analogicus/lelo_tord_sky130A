*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bias_1p2u_lpe.spi
#else
.include ../../../work/xsch/bias_1p2u.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.csparam voltage_supply_csparam = {vdda}

.param delay = 10ns
.param rise = 1ns
.param width = 100ns
.param fall = 1ns

.param sleep_signal = 0V
.csparam sleep_signal_csparam = {sleep_signal}

.param simulation_length = 50ns
.csparam simulation_length_csparam = {simulation_length}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0 dc 0V
VDD VDD VSS dc {AVDD}
VSLEEP SLEEP VSS dc {sleep_signal}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

set sim_len = {$&simulation_length_csparam}
set slp_sig = {$&sleep_signal_csparam}
set vsup = {$&voltage_supply_csparam}

optran 0 0 0 1ns 1us 0
tran 1ns $sim_len 10ps
write 

alterparam sleep_signal = {$vsup}
reset

optran 0 0 0 1ns 1us 0
tran 1ns $sim_len 10ps
write {cicname}_sleep_high.raw

quit

.endc

.end
