*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_tmp_core_and_cmp_lpe.spi
#else
.include ../../../work/xsch/TB_tmp_core_and_cmp.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS     VSS    0   dc 0V
VDD     VDD    VSS dc {AVDD}
VSLEEP  SLEEP  VSS dc 0V
IPTAT   IPTAT  VSS dc 1uA
VRST    RST    VSS pwl 0s 0V 900ns 0V 910ns {AVDD} 920ns 0V
VREF    REF    VSS dc 1V
VCMP_P1 CMP_P1 VSS dc {AVDD}
VCMP_P2 CMP_P2 VSS dc 0V

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.option savecurrents
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 10n 10p
write
quit


.endc

.end
